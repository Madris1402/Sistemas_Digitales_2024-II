// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Wed Mar 13 17:53:26 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module contador_cuatro_bits (
    reset,clock,
    output1,output2,output3,output4);

    input reset;
    input clock;
    tri0 reset;
    output output1;
    output output2;
    output output3;
    output output4;
    reg output1;
    reg output2;
    reg output3;
    reg output4;
    reg [15:0] fstate;
    reg [15:0] reg_fstate;
    parameter state5=0,state14=1,state10=2,state9=3,state1=4,state3=5,state8=6,state7=7,state4=8,state6=9,state11=10,state12=11,state13=12,state16=13,state2=14,state15=15;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset)
    begin
        if (reset) begin
            reg_fstate <= state1;
            output1 <= 1'b0;
            output2 <= 1'b0;
            output3 <= 1'b0;
            output4 <= 1'b0;
        end
        else begin
            output1 <= 1'b0;
            output2 <= 1'b0;
            output3 <= 1'b0;
            output4 <= 1'b0;
            case (fstate)
                state5: begin
                    reg_fstate <= state6;

                    output4 <= 1'b0;

                    output2 <= 1'b1;

                    output3 <= 1'b0;

                    output1 <= 1'b0;
                end
                state14: begin
                    reg_fstate <= state15;

                    output4 <= 1'b1;

                    output2 <= 1'b1;

                    output3 <= 1'b0;

                    output1 <= 1'b1;
                end
                state10: begin
                    reg_fstate <= state11;

                    output4 <= 1'b1;

                    output2 <= 1'b0;

                    output3 <= 1'b0;

                    output1 <= 1'b1;
                end
                state9: begin
                    reg_fstate <= state10;

                    output4 <= 1'b0;

                    output2 <= 1'b0;

                    output3 <= 1'b0;

                    output1 <= 1'b1;
                end
                state1: begin
                    reg_fstate <= state2;

                    output4 <= 1'b0;

                    output2 <= 1'b0;

                    output3 <= 1'b0;

                    output1 <= 1'b0;
                end
                state3: begin
                    reg_fstate <= state4;

                    output4 <= 1'b0;

                    output2 <= 1'b0;

                    output3 <= 1'b1;

                    output1 <= 1'b0;
                end
                state8: begin
                    reg_fstate <= state9;

                    output4 <= 1'b1;

                    output2 <= 1'b1;

                    output3 <= 1'b1;

                    output1 <= 1'b0;
                end
                state7: begin
                    reg_fstate <= state8;

                    output4 <= 1'b0;

                    output2 <= 1'b1;

                    output3 <= 1'b1;

                    output1 <= 1'b0;
                end
                state4: begin
                    reg_fstate <= state5;

                    output4 <= 1'b1;

                    output2 <= 1'b0;

                    output3 <= 1'b1;

                    output1 <= 1'b0;
                end
                state6: begin
                    reg_fstate <= state7;

                    output4 <= 1'b1;

                    output2 <= 1'b1;

                    output3 <= 1'b0;

                    output1 <= 1'b0;
                end
                state11: begin
                    reg_fstate <= state12;

                    output1 <= 1'b1;
                    output1 <= 1'b0;
                    output1 <= 1'b1;
                    output1 <= 1'b0;
                end
                state12: begin
                    reg_fstate <= state13;

                    output4 <= 1'b1;

                    output2 <= 1'b0;

                    output3 <= 1'b1;

                    output1 <= 1'b1;
                end
                state13: begin
                    reg_fstate <= state14;

                    output4 <= 1'b0;

                    output2 <= 1'b1;

                    output3 <= 1'b0;

                    output1 <= 1'b1;
                end
                state16: begin
                    reg_fstate <= state1;

                    output4 <= 1'b1;

                    output2 <= 1'b1;

                    output3 <= 1'b1;

                    output1 <= 1'b1;
                end
                state2: begin
                    reg_fstate <= state3;

                    output4 <= 1'b1;

                    output2 <= 1'b0;

                    output3 <= 1'b0;

                    output1 <= 1'b0;
                end
                state15: begin
                    reg_fstate <= state16;

                    output4 <= 1'b0;

                    output2 <= 1'b1;

                    output3 <= 1'b1;

                    output1 <= 1'b1;
                end
                default: begin
                    output1 <= 1'bx;
                    output2 <= 1'bx;
                    output3 <= 1'bx;
                    output4 <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // contador_cuatro_bits
