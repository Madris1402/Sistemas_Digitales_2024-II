library verilog;
use verilog.vl_types.all;
entity flipflopJK_negedge1_vlg_vec_tst is
end flipflopJK_negedge1_vlg_vec_tst;
