library verilog;
use verilog.vl_types.all;
entity divisor_vlg_check_tst is
    port(
        ckd             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end divisor_vlg_check_tst;
