library verilog;
use verilog.vl_types.all;
entity compuerta_and_vlg_vec_tst is
end compuerta_and_vlg_vec_tst;
