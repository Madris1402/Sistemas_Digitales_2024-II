library verilog;
use verilog.vl_types.all;
entity contador_cuatro_bits_vlg_vec_tst is
end contador_cuatro_bits_vlg_vec_tst;
