library verilog;
use verilog.vl_types.all;
entity flipflopJK_negedge1_vlg_check_tst is
    port(
        CLK2            : in     vl_logic;
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end flipflopJK_negedge1_vlg_check_tst;
