library verilog;
use verilog.vl_types.all;
entity flipflop_JK_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        J               : in     vl_logic;
        K               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end flipflop_JK_vlg_sample_tst;
