library verilog;
use verilog.vl_types.all;
entity tbt_vlg_check_tst is
    port(
        ckd             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end tbt_vlg_check_tst;
