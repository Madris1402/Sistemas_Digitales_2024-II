library verilog;
use verilog.vl_types.all;
entity latch_D_vlg_vec_tst is
end latch_D_vlg_vec_tst;
