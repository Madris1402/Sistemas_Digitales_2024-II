library verilog;
use verilog.vl_types.all;
entity latch_RS_nandEN_vlg_vec_tst is
end latch_RS_nandEN_vlg_vec_tst;
