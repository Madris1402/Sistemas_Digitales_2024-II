library verilog;
use verilog.vl_types.all;
entity latches_vlg_vec_tst is
end latches_vlg_vec_tst;
