library verilog;
use verilog.vl_types.all;
entity tbt_vlg_vec_tst is
end tbt_vlg_vec_tst;
