// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Fri Mar 15 00:28:26 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module contador_cuatro_bits (
    reset,clock,input1,
    output1,output2,output3,output4);

    input reset;
    input clock;
    input input1;
    tri0 reset;
    tri0 input1;
    output output1;
    output output2;
    output output3;
    output output4;
    reg output1;
    reg output2;
    reg output3;
    reg output4;
    reg [15:0] fstate;
    reg [15:0] reg_fstate;
    parameter state16=0,state15=1,state3=2,state14=3,state4=4,state13=5,state12=6,state5=7,state11=8,state10=9,state7=10,state8=11,state1=12,state2=13,state9=14,state6=15;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or input1)
    begin
        if (reset) begin
            reg_fstate <= state1;
            output1 <= 1'b0;
            output2 <= 1'b0;
            output3 <= 1'b0;
            output4 <= 1'b0;
        end
        else begin
            output1 <= 1'b0;
            output2 <= 1'b0;
            output3 <= 1'b0;
            output4 <= 1'b0;
            case (fstate)
                state16: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state1;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state15;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state16;

                    output4 <= 1'b1;

                    output3 <= 1'b1;

                    output2 <= 1'b1;

                    output1 <= 1'b1;
                end
                state15: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state16;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state14;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state15;

                    output4 <= 1'b0;

                    output3 <= 1'b1;

                    output2 <= 1'b1;

                    output1 <= 1'b1;
                end
                state3: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state4;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    output4 <= 1'b0;

                    output3 <= 1'b1;

                    output2 <= 1'b0;

                    output1 <= 1'b0;
                end
                state14: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state15;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state13;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state14;

                    output4 <= 1'b1;

                    output3 <= 1'b0;

                    output2 <= 1'b1;

                    output1 <= 1'b1;
                end
                state4: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state5;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    output4 <= 1'b1;

                    output3 <= 1'b1;

                    output2 <= 1'b0;

                    output1 <= 1'b0;
                end
                state13: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state12;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state14;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state13;

                    output4 <= 1'b0;

                    output3 <= 1'b0;

                    output2 <= 1'b1;

                    output1 <= 1'b1;
                end
                state12: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state13;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state11;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state12;

                    output4 <= 1'b1;

                    output3 <= 1'b1;

                    output2 <= 1'b0;

                    output1 <= 1'b1;
                end
                state5: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state4;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    output4 <= 1'b0;

                    output3 <= 1'b0;

                    output2 <= 1'b1;

                    output1 <= 1'b0;
                end
                state11: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state12;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state10;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state11;

                    output4 <= 1'b0;

                    output3 <= 1'b1;

                    output2 <= 1'b0;

                    output1 <= 1'b1;
                end
                state10: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state9;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state11;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state10;

                    output4 <= 1'b1;

                    output3 <= 1'b0;

                    output2 <= 1'b0;

                    output1 <= 1'b1;
                end
                state7: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state8;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state7;

                    output4 <= 1'b0;

                    output3 <= 1'b1;

                    output2 <= 1'b1;

                    output1 <= 1'b0;
                end
                state8: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state7;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state9;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state8;

                    output4 <= 1'b1;

                    output3 <= 1'b1;

                    output2 <= 1'b1;

                    output1 <= 1'b0;
                end
                state1: begin
                    if ((input1 == 1'b0))
                        reg_fstate <= state16;
                    else if ((input1 == 1'b1))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    output4 <= 1'b0;

                    output3 <= 1'b0;

                    output2 <= 1'b0;

                    output1 <= 1'b0;
                end
                state2: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state3;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    output4 <= 1'b1;

                    output3 <= 1'b0;

                    output2 <= 1'b0;

                    output1 <= 1'b0;
                end
                state9: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state10;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state8;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state9;

                    output4 <= 1'b0;

                    output3 <= 1'b0;

                    output2 <= 1'b0;

                    output1 <= 1'b1;
                end
                state6: begin
                    if ((input1 == 1'b1))
                        reg_fstate <= state7;
                    else if ((input1 == 1'b0))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state6;

                    output4 <= 1'b1;

                    output3 <= 1'b0;

                    output2 <= 1'b1;

                    output1 <= 1'b0;
                end
                default: begin
                    output1 <= 1'bx;
                    output2 <= 1'bx;
                    output3 <= 1'bx;
                    output4 <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // contador_cuatro_bits
