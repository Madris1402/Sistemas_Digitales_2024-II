library verilog;
use verilog.vl_types.all;
entity lsr_vlg_vec_tst is
end lsr_vlg_vec_tst;
