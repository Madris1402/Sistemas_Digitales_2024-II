library verilog;
use verilog.vl_types.all;
entity seqdiv_vlg_sample_tst is
    port(
        ck              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end seqdiv_vlg_sample_tst;
