library verilog;
use verilog.vl_types.all;
entity compuerta_and_vlg_check_tst is
    port(
        s1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end compuerta_and_vlg_check_tst;
