library verilog;
use verilog.vl_types.all;
entity SM2_vlg_vec_tst is
end SM2_vlg_vec_tst;
