library verilog;
use verilog.vl_types.all;
entity flipflopJK_negedge1 is
    port(
        CLK2            : out    vl_logic;
        CLK             : in     vl_logic;
        E1              : in     vl_logic;
        Q               : out    vl_logic
    );
end flipflopJK_negedge1;
