library verilog;
use verilog.vl_types.all;
entity flipflop_D_vlg_vec_tst is
end flipflop_D_vlg_vec_tst;
