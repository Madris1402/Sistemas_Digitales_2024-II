library verilog;
use verilog.vl_types.all;
entity flipflop_d_vlg_vec_tst is
end flipflop_d_vlg_vec_tst;
