library verilog;
use verilog.vl_types.all;
entity Pastillero_vlg_vec_tst is
end Pastillero_vlg_vec_tst;
