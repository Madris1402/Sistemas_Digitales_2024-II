library verilog;
use verilog.vl_types.all;
entity compuerta_and_vlg_sample_tst is
    port(
        e1              : in     vl_logic;
        e2              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end compuerta_and_vlg_sample_tst;
