library verilog;
use verilog.vl_types.all;
entity rx_vlg_vec_tst is
end rx_vlg_vec_tst;
