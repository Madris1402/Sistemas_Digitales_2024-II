library verilog;
use verilog.vl_types.all;
entity divisor_vlg_sample_tst is
    port(
        ck              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end divisor_vlg_sample_tst;
