library verilog;
use verilog.vl_types.all;
entity cascada_JK_vlg_vec_tst is
end cascada_JK_vlg_vec_tst;
