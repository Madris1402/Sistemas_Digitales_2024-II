library verilog;
use verilog.vl_types.all;
entity prot_vlg_vec_tst is
end prot_vlg_vec_tst;
