library verilog;
use verilog.vl_types.all;
entity flipflop_T_vlg_vec_tst is
end flipflop_T_vlg_vec_tst;
