library verilog;
use verilog.vl_types.all;
entity compuerta_and is
    port(
        e1              : in     vl_logic;
        e2              : in     vl_logic;
        s1              : out    vl_logic
    );
end compuerta_and;
