library verilog;
use verilog.vl_types.all;
entity latch_JK_vlg_vec_tst is
end latch_JK_vlg_vec_tst;
