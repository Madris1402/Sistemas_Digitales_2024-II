library verilog;
use verilog.vl_types.all;
entity seqdiv_vlg_vec_tst is
end seqdiv_vlg_vec_tst;
