library verilog;
use verilog.vl_types.all;
entity flipflop_RS_nor_vlg_vec_tst is
end flipflop_RS_nor_vlg_vec_tst;
