library verilog;
use verilog.vl_types.all;
entity flipflop_JK_vlg_vec_tst is
end flipflop_JK_vlg_vec_tst;
